version https://git-lfs.github.com/spec/v1
oid sha256:26f4cb0fab3819a8a4de2c5c6bf46eb47da8115440c0e43868be58b949afa244
size 429968
