version https://git-lfs.github.com/spec/v1
oid sha256:b18b2ff9d7ce5f411c65ac76a0338350e6956840d1f5df729210b39b541ad63f
size 568853
