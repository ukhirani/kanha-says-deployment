version https://git-lfs.github.com/spec/v1
oid sha256:1edc00c4f4e40fc076fb38cadace7d9b8e431658ef7a9fe5c9f2da1af02231f4
size 562271
