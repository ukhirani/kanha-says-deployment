version https://git-lfs.github.com/spec/v1
oid sha256:334503d01e43313b5749dd81cedb91b0820217f40b13699ed8bf0320dfe56be6
size 317764
