version https://git-lfs.github.com/spec/v1
oid sha256:4d9a350ad15f72c1b825d57d6d4eb6fb5a22230b51a88aec53472cb355a2d829
size 336578
