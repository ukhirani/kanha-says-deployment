version https://git-lfs.github.com/spec/v1
oid sha256:94e8a2072fa4ca5e078b1ef887f5a4f1f5fd41be6be240613a91a0c3c9b93fbb
size 74752
