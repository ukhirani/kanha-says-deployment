version https://git-lfs.github.com/spec/v1
oid sha256:661ebd2799d09eb5a6f65e6639383313fc47579399e76977830427b34f758160
size 147626
