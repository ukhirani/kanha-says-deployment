version https://git-lfs.github.com/spec/v1
oid sha256:4094bdd5d2286c4d185c51d9381497b24f6010a128a987a9e7c476d0d9d94252
size 586195
