version https://git-lfs.github.com/spec/v1
oid sha256:3ab201c1d70b2c9ec35592479ea83275eaba1fca9e84cd1af151f4bdbfd4a10a
size 150668
