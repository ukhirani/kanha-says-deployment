version https://git-lfs.github.com/spec/v1
oid sha256:787ca5db33c87a528e9f130cecc0da162571cfd5d14fa46f63cbb5c8eae89144
size 176798
